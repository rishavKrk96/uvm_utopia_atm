// Code your design here
`include "squat.sv"
`include "utopia1_atm_rx.sv"
`include "utopia1_atm_tx.sv"