// Code your testbench here
// or browse Examples
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "definitions.sv"  // include external definitions
`include "config.svh"
`include "utopia.sv"
`include "top.sv"
`include "cpu_ifc.sv"
`include "LookupTable.sv"
`include "atm_cell.sv"
`include "sequence.svh"
`include "driver.svh"
`include "monitor.svh"
`include "sequencer.svh"
`include "cpu_ifc.sv"
`include "cpu_driver.svh"
`include "agent.svh"
`include "scoreboard.svh"
`include "coverage.svh"
`include "environment.svh"
`include "test.sv"


